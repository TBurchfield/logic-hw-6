module hw6_tb(
);

endmodule
